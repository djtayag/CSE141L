package Definitions;

   typedef enum logic [3:0] {
       ADD,
       LSH,
       RSH,
       XOR,
       AND,
       SUB,
       CLR
   } op_mne;

endpackage // Definitions
